module NOT(input[7:0] inA, output[7:0] out);
    assign out = ~inA;
endmodule