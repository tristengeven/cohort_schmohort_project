// logic op not
module NOT(input[15:0] inA, output[15:0] out);
    assign out = ~inA; // not
endmodule