module XOR(input[7:0] inA, inB, output[7:0] out);
    assign out = inA ^ inB;
endmodule