// logic op xor
module XOR(input[15:0] A, B, output[15:0] out);
    assign out = A ^ B; // xor
endmodule