// logic op xor
module XOR(input[15:0] inA, inB, output[15:0] out);
    assign out = inA ^ inB; // xor
endmodule