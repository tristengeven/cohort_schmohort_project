// logic op not
module NOT(input[15:0] A, output[15:0] out);
    assign out = ~A; // not
endmodule